
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/BreakWhile/top.sv:1.1-10.10" *)
module top(a);
  (* src = "/root/synlig/synlig/tests/simple_tests/BreakWhile/top.sv:1.23-1.24" *)
  output [31:0] a;
  wire [31:0] a;
  assign a = 32'd128;
endmodule
