
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/FunctionCallsFunctionWithIndexedPartSelectAsArgument/top.sv:13.1-15.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/FunctionCallsFunctionWithIndexedPartSelectAsArgument/top.sv:13.32-13.33" *)
  output [15:0] o;
  wire [15:0] o;
  assign o = 16'hxxcd;
endmodule
