
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypedefInModulePort/top.sv:6.1-8.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefInModulePort/top.sv:6.32-6.33" *)
  (* wiretype = "\\word" *)
  output [7:0] o;
  wire [7:0] o;
  assign o = 8'h5c;
endmodule
