
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/event_implicit_expression_list/event_implicit.sv:6.1-14.10" *)
module top();
  (* src = "/root/synlig/synlig/tests/simple_tests/event_implicit_expression_list/event_implicit.sv:7.7-7.8" *)
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/event_implicit_expression_list/event_implicit.sv:8.7-8.8" *)
  wire b;
  (* src = "/root/synlig/synlig/tests/simple_tests/event_implicit_expression_list/event_implicit.sv:9.7-9.8" *)
  wire c;
  (* src = "/root/synlig/synlig/tests/simple_tests/event_implicit_expression_list/event_implicit.sv:10.7-10.8" *)
  wire d;
  (* src = "/root/synlig/synlig/tests/simple_tests/event_implicit_expression_list/event_implicit.sv:11.6-11.9" *)
  wire out;
  assign a = 1'h0;
  assign b = 1'h0;
  assign c = 1'h0;
  assign d = 1'h0;
  assign out = 1'h0;
endmodule
