
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/BitsCallOnParametetrizedTypeFromPackage/top.sv:6.1-10.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/BitsCallOnParametetrizedTypeFromPackage/top.sv:6.23-6.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd10;
endmodule
