
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ImportFunction/top.sv:12.1-14.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ImportFunction/top.sv:12.23-12.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd5;
endmodule
