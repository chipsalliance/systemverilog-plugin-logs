
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumFirst/top.sv:1.1-6.10" *)
module top(o);
  (* enum_value_00000000000000000000000000000001 = "\\a" *)
  (* enum_value_00000000000000000000000000000010 = "\\b" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumFirst/top.sv:4.12-4.13" *)
  (* wiretype = "\\my_enum" *)
  wire [31:0] e;
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumFirst/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign e = o;
endmodule
