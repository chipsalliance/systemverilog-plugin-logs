
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CastClog2/top.sv:1.1-6.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CastClog2/top.sv:1.31-1.32" *)
  output [1:0] o;
  wire [1:0] o;
  assign o = 2'h3;
endmodule
