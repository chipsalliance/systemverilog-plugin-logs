
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EmptyTask/top.sv:6.1-11.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/EmptyTask/top.sv:6.19-6.20" *)
  output o;
  wire o;
  assign o = 1'h1;
endmodule
