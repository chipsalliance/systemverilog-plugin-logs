
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ParameterPackedArraySurelogSubstitution/top.sv:3.1-7.10" *)
module top(a);
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterPackedArraySurelogSubstitution/top.sv:3.30-3.31" *)
  output [3:0] a;
  wire [3:0] a;
  assign a = 4'h1;
endmodule
