
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/MultiAssignmentPatternOfConcat/top.sv:1.1-6.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/MultiAssignmentPatternOfConcat/top.sv:4.8-4.9" *)
  wire [191:0] n;
  (* src = "/root/synlig/synlig/tests/simple_tests/MultiAssignmentPatternOfConcat/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign n = 192'h000000040000000500000004000000050000000400000005;
  assign o = 32'd4;
endmodule
