
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/DeclarationInFor/top.sv:1.1-12.16" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/DeclarationInFor/top.sv:1.25-1.26" *)
  output o;
  wire o;
  assign o = 1'h1;
endmodule
