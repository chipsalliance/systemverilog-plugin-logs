
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/simple_unary_op_plus/simple_unary_op_plus.sv:6.1-8.10" *)
module top(a, b);
  (* src = "/root/synlig/synlig/tests/simple_tests/simple_unary_op_plus/simple_unary_op_plus.sv:6.24-6.25" *)
  input [3:0] a;
  wire [3:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/simple_unary_op_plus/simple_unary_op_plus.sv:6.40-6.41" *)
  output [3:0] b;
  wire [3:0] b;
  assign b = a;
endmodule
