
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/Function2Returns/top.sv:8.1-10.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/Function2Returns/top.sv:8.19-8.20" *)
  output o;
  wire o;
  assign o = 1'h1;
endmodule
