
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumInGenblock/top.sv:1.1-31.10" *)
module top();
endmodule
