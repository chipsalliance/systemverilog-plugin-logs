
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/PackedInGenblock/top.sv:6.1-12.10" *)
module top();
endmodule
