
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/AnonStructs/top.sv:1.1-18.10" *)
module top(b);
  (* src = "/root/synlig/synlig/tests/simple_tests/AnonStructs/top.sv:0.0-0.0" *)
  (* wiretype = "\\a" *)
  wire [3:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/AnonStructs/top.sv:1.25-1.26" *)
  output [3:0] b;
  wire [3:0] b;
  assign a = 4'h5;
  assign b = 4'h5;
endmodule
