
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypedefedRangedFunctionReturn/top.sv:1.1-8.10" *)
module top(a, b);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefedRangedFunctionReturn/top.sv:1.32-1.33" *)
  output [31:0] a;
  wire [31:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefedRangedFunctionReturn/top.sv:1.35-1.36" *)
  output [31:0] b;
  wire [31:0] b;
  assign a = 32'd0;
  assign b = 32'd1;
endmodule
