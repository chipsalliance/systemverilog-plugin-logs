
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/unary_op_plus/unary_op_plus.sv:6.1-12.10" *)
module top();
  (* src = "/root/synlig/synlig/tests/simple_tests/unary_op_plus/unary_op_plus.sv:7.5-7.11" *)
  wire [31:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/unary_op_plus/unary_op_plus.sv:8.5-8.10" *)
  wire [31:0] b;
  assign a = 32'd5;
  assign b = 32'd5;
endmodule
