
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TaskExportDPI/top.sv:1.1-12.10" *)
module top(a);
  (* src = "/root/synlig/synlig/tests/simple_tests/TaskExportDPI/top.sv:1.23-1.24" *)
  output [31:0] a;
  wire [31:0] a;
  (* nosync = 32'd1 *)
  (* src = "/root/synlig/synlig/tests/simple_tests/TaskExportDPI/top.sv:7.49-7.50" *)
  wire [31:0] \get_2$func$/root/synlig/synlig/tests/simple_tests/TaskExportDPI/top.sv:10$1.x ;
  assign \get_2$func$/root/synlig/synlig/tests/simple_tests/TaskExportDPI/top.sv:10$1.x  = a;
endmodule
