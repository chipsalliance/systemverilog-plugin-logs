
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/AnonymousUnion/top.sv:1.1-11.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/AnonymousUnion/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  (* src = "/root/synlig/synlig/tests/simple_tests/AnonymousUnion/top.sv:0.0-0.0" *)
  (* wiretype = "\\un" *)
  wire [31:0] un;
  assign o = 32'd1;
  assign un = 32'd1;
endmodule
