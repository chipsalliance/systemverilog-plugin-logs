
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/PatternStruct/top.sv:1.1-7.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/PatternStruct/top.sv:1.31-1.32" *)
  output [7:0] o;
  wire [7:0] o;
  (* src = "/root/synlig/synlig/tests/simple_tests/PatternStruct/top.sv:5.14-5.15" *)
  (* wiretype = "\\my_struct" *)
  wire [7:0] s;
  assign o = 8'h7d;
  assign s = 8'h7d;
endmodule
