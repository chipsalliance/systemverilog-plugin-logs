
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/BitsCallOnVar/top.sv:1.1-9.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/BitsCallOnVar/top.sv:6.29-6.44" *)
  wire [31:0] dr_q;
  (* src = "/root/synlig/synlig/tests/simple_tests/BitsCallOnVar/top.sv:1.32-1.33" *)
  output [31:0] o;
  wire [31:0] o;
  assign dr_q = 32'd43981;
  assign o = 32'd43981;
endmodule
