
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CastExpression/top.sv:1.1-8.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CastExpression/top.sv:4.17-4.27" *)
  wire [15:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/CastExpression/top.sv:1.31-1.32" *)
  output [4:0] o;
  wire [4:0] o;
  assign a = 16'h00ab;
  assign o = 5'h0b;
endmodule
