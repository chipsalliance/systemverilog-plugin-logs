
(* cells_not_processed =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/FileLevelParameter/top.sv:2.1-8.10" *)
module top();
  reg \$auto$verilog_backend.cc:2352:dump_module$3  = 0;
  always @* begin
    if (\$auto$verilog_backend.cc:2352:dump_module$3 ) begin end
    (* src = "/root/synlig/synlig/tests/simple_tests/FileLevelParameter/top.sv:4.5-6.8" *)
        end
  end
  always @* begin
  end
endmodule
