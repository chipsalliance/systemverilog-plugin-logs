
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/2DeclarationsInFor/top.sv:1.1-13.16" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/2DeclarationsInFor/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd3;
endmodule
