
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumConcat/dut.v:7.1-19.10" *)
module dut(a0);
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumConcat/dut.v:7.12-7.14" *)
  input a0;
  wire a0;
endmodule
