
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/BitsCallOnSubArray/top.sv:10.1-13.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/BitsCallOnSubArray/top.sv:10.23-10.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd16;
endmodule
