
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/BindModuleWithInputPortsInGenScope/top.sv:7.1-12.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/BindModuleWithInputPortsInGenScope/top.sv:7.23-7.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd10;
endmodule
