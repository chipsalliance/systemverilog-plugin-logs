
(* src = "/root/synlig/synlig/tests/simple_tests/ImportedEnumCast/top.sv:13.5-15.23" *)
module \$paramod\generic_flop\ResetValue=4'1001 ();
endmodule

(* src = "/root/synlig/synlig/tests/simple_tests/ImportedEnumCast/top.sv:21.3-23.19" *)
module \$paramod\prim_flop\ResetValue=4'1001 ();
endmodule

(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ImportedEnumCast/top.sv:18.1-25.10" *)
module top();
endmodule
