
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/UnpackedArray/top.sv:1.1-5.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/UnpackedArray/top.sv:1.23-1.24" *)
  output [383:0] o;
  wire [383:0] o;
  assign o = 384'h000000000000000100000002000000030000000a0000000b0000000c0000000d00000014000000150000001600000017;
endmodule
