
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/StructPackedArray/top.sv:1.1-8.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/StructPackedArray/top.sv:6.23-6.43" *)
  (* wiretype = "\\filter_ctl_t" *)
  wire [19:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/StructPackedArray/top.sv:1.31-1.32" *)
  output [9:0] o;
  wire [9:0] o;
  assign a = 20'h03c00;
  assign o = 10'h00f;
endmodule
