
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ImportTypeOfPort/top.sv:6.1-10.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ImportTypeOfPort/top.sv:7.19-7.20" *)
  (* wiretype = "\\lc_tx_t" *)
  output [3:0] o;
  wire [3:0] o;
  assign o = 4'h5;
endmodule
