
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ReferencedPackageParameterInEnum/top.sv:11.1-13.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ReferencedPackageParameterInEnum/top.sv:11.23-11.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd24;
endmodule
