
(* src = "/root/synlig/synlig/tests/simple_tests/EnumItemReimport/top.sv:15.3-15.10" *)
module M();
endmodule

(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumItemReimport/top.sv:14.1-16.10" *)
module top();
endmodule
