
(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnum/top.sv:25.3-29.5" *)
module \$paramod$808d8cab74cca023878377ed823b6ee10422a46f\test_module (state_i);
  (* enum_value_100100001 = "\\enum_bar_e$enum3.\\BarVariant" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnum/top.sv:4.24-4.31" *)
  (* wiretype = "\\enum_bar_e" *)
  input [8:0] state_i;
  wire [8:0] state_i;
endmodule

(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnum/top.sv:14.3-18.5" *)
module \$paramod$ae563f53012966872350ccb3ebfb43ff1886ac87\test_module (state_i);
  (* enum_value_10010101 = "\\enum_foo_e$enum2.\\FooVariant" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnum/top.sv:4.24-4.31" *)
  (* wiretype = "\\enum_foo_e" *)
  input [7:0] state_i;
  wire [7:0] state_i;
endmodule

(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnum/top.sv:8.1-30.10" *)
module top();
endmodule
