
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CastLogic/top.sv:1.1-3.10" *)
module top(clk, o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CastLogic/top.sv:1.18-1.21" *)
  input clk;
  wire clk;
  (* src = "/root/synlig/synlig/tests/simple_tests/CastLogic/top.sv:1.36-1.37" *)
  output o;
  wire o;
  assign o = 1'h1;
endmodule
