
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumArray/top.sv:7.1-10.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumArray/top.sv:7.23-7.24" *)
  output [31:0] o;
  wire [31:0] o;
  (* enum_value_1010 = "\\On" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumArray/top.sv:8.26-8.46" *)
  (* wiretype = "\\lc_tx_t" *)
  wire [31:0] x;
  assign o = 32'd2863311530;
  assign x = 32'd2863311530;
endmodule
