
(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnumOfParametrizedWidth/top.sv:18.3-22.5" *)
module \$paramod$b2778081825e52137dcae6c464d171bf273c42c0\test_module (state_i);
  (* enum_value_100100001 = "\\state_e$enum1.\\StActive" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnumOfParametrizedWidth/top.sv:4.24-4.31" *)
  (* wiretype = "\\state_e" *)
  input [8:0] state_i;
  wire [8:0] state_i;
endmodule

(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithEnumOfParametrizedWidth/top.sv:8.1-24.16" *)
module top();
endmodule
