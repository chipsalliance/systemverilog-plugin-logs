
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumVariantInPackage/top.sv:14.1-16.10" *)
module top(i, o);
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumVariantInPackage/top.sv:14.24-14.25" *)
  input i;
  wire i;
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumVariantInPackage/top.sv:14.40-14.41" *)
  output o;
  wire o;
  (* enum_value_0 = "\\Off" *)
  (* enum_value_1 = "\\On" *)
  (* nosync = 32'd1 *)
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumVariantInPackage/top.sv:8.46-8.49" *)
  (* wiretype = "\\lc_tx_t" *)
  wire \test_package::test_true$func$/root/synlig/synlig/tests/simple_tests/EnumVariantInPackage/top.sv:15$2.val ;
  assign o = i;
  assign \test_package::test_true$func$/root/synlig/synlig/tests/simple_tests/EnumVariantInPackage/top.sv:15$2.val  = 1'hx;
endmodule
