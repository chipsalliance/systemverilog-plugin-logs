
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/GenIfInside/top.sv:13.1-33.10" *)
module top(out);
  (* src = "/root/synlig/synlig/tests/simple_tests/GenIfInside/top.sv:18.16-18.19" *)
  output [31:0] out;
  wire [31:0] out;
  assign out = 32'd0;
endmodule
