
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ScopeOverwriting/top.sv:1.1-18.10" *)
module top();
endmodule
