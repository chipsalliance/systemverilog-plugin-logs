
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/BitSelect2ndBitOfPattern/top.sv:1.1-4.10" *)
module top(a);
  (* src = "/root/synlig/synlig/tests/simple_tests/BitSelect2ndBitOfPattern/top.sv:1.25-1.26" *)
  output a;
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/BitSelect2ndBitOfPattern/top.sv:2.10-2.11" *)
  wire [1:0] x;
  assign a = 1'h1;
  assign x = 2'h2;
endmodule
