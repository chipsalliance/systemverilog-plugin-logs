
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/VarInFor/top.sv:12.1-14.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/VarInFor/top.sv:12.27-12.28" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd3;
endmodule
