
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CastToSumOfConstants/top.sv:1.1-5.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CastToSumOfConstants/top.sv:1.31-1.32" *)
  output [2:0] o;
  wire [2:0] o;
  assign o = 3'h7;
endmodule
