
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/Longint/top.sv:1.1-3.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/Longint/top.sv:1.27-1.28" *)
  output [63:0] o;
  wire [63:0] o;
  assign o = 64'h0000000000000001;
endmodule
