
(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithLogic/top.sv:21.3-25.5" *)
module \$paramod$71a5c9f5858ab9c319d21440db8ec918fe727532\test_module (state_i);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithLogic/top.sv:4.24-4.31" *)
  (* wiretype = "\\foo_type" *)
  input [2:0] state_i;
  wire [2:0] state_i;
endmodule

(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithLogic/top.sv:12.3-16.5" *)
module \$paramod$b2778081825e52137dcae6c464d171bf273c42c0\test_module (state_i);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithLogic/top.sv:4.24-4.31" *)
  (* wiretype = "\\state_e" *)
  input state_i;
  wire state_i;
endmodule

(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypeParameterAsPortTypeWithLogic/top.sv:8.1-32.10" *)
module top();
endmodule
