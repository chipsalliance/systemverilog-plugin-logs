
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypedefStructArray/top.sv:1.1-7.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefStructArray/top.sv:5.19-5.20" *)
  (* wiretype = "\\struct_array_t" *)
  wire [31:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefStructArray/top.sv:1.32-1.33" *)
  output [31:0] o;
  wire [31:0] o;
  assign a = 32'd4294967295;
  assign o = 32'd4294967295;
endmodule
