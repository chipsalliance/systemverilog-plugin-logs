
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumConcatenatedConst/top.sv:10.1-12.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumConcatenatedConst/top.sv:10.32-10.33" *)
  output [63:0] o;
  wire [63:0] o;
  assign o = 64'h0000000100000001;
endmodule
