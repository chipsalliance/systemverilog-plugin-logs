
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypedefAliasInPackage/top.sv:10.1-15.10" *)
module top(o);
  (* enum_value_1010 = "\\On" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefAliasInPackage/top.sv:11.25-11.50" *)
  (* wiretype = "\\lc_tx_e" *)
  wire [3:0] lc_en_i;
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefAliasInPackage/top.sv:10.31-10.32" *)
  output [3:0] o;
  wire [3:0] o;
  assign lc_en_i = 4'ha;
  assign o = 4'ha;
endmodule
