
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/StructParameterInitializedWithPatternAndReferenced/top.sv:13.1-15.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/StructParameterInitializedWithPatternAndReferenced/top.sv:13.23-13.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd3;
endmodule
