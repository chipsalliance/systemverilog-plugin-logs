
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ConstSizes/dut.v:1.1-6.10" *)
module dut(a, b, c, d);
  (* src = "/root/synlig/synlig/tests/simple_tests/ConstSizes/dut.v:1.32-1.33" *)
  output [63:0] a;
  wire [63:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/ConstSizes/dut.v:1.54-1.55" *)
  output [63:0] b;
  wire [63:0] b;
  (* src = "/root/synlig/synlig/tests/simple_tests/ConstSizes/dut.v:1.76-1.77" *)
  output [63:0] c;
  wire [63:0] c;
  (* src = "/root/synlig/synlig/tests/simple_tests/ConstSizes/dut.v:1.98-1.99" *)
  output [63:0] d;
  wire [63:0] d;
  assign a = 64'h6ad5d6150952103c;
  assign b = 64'h6ad5d6150952103c;
  assign c = 64'hadb52acaaaaaaaae;
  assign d = 64'hacbf74cfa4b5a09b;
endmodule
