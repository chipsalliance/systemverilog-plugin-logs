
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/AssignSumOfConstants/top.sv:1.1-3.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/AssignSumOfConstants/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd3;
endmodule
