
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CastStructArray/top.sv:1.1-12.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CastStructArray/top.sv:8.17-8.27" *)
  wire [15:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/CastStructArray/top.sv:1.31-1.32" *)
  output [5:0] o;
  wire [5:0] o;
  assign a = 16'h00ab;
  assign o = 6'h2b;
endmodule
