
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypedefedFunctionReturn/top.sv:1.1-8.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefedFunctionReturn/top.sv:1.32-1.33" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd43981;
endmodule
