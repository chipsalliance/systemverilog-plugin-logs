
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.1-28.10" *)
module top(a, b, c, d, e, f, g, h, i, j, k, l);
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.25-1.26" *)
  output a;
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.28-1.29" *)
  output b;
  wire b;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.31-1.32" *)
  output c;
  wire c;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.34-1.35" *)
  output d;
  wire d;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.37-1.38" *)
  output e;
  wire e;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.40-1.41" *)
  output f;
  wire f;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.43-1.44" *)
  output g;
  wire g;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.46-1.47" *)
  output h;
  wire h;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.49-1.50" *)
  output i;
  wire i;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.52-1.53" *)
  output j;
  wire j;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.55-1.56" *)
  output k;
  wire k;
  (* src = "/root/synlig/synlig/tests/simple_tests/compound_assignments/top.sv:1.58-1.59" *)
  output l;
  wire l;
  assign a = 1'h0;
  assign b = 1'h0;
  assign c = 1'h1;
  assign d = 1'h0;
  assign e = 1'h0;
  assign f = 1'h0;
  assign g = 1'h0;
  assign h = 1'h1;
  assign i = 1'h0;
  assign j = 1'h1;
  assign k = 1'h0;
  assign l = 1'h0;
endmodule
