
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/GenblockPackedAccess/top.sv:1.1-13.10" *)
module top();
  (* src = "/root/synlig/synlig/tests/simple_tests/GenblockPackedAccess/top.sv:11.11-11.12" *)
  wire \n.x.foo.a ;
  (* src = "/root/synlig/synlig/tests/simple_tests/GenblockPackedAccess/top.sv:12.11-12.12" *)
  wire \n.x.foo.b ;
  assign \n.x.foo.a  = 1'h0;
  assign \n.x.foo.b  = 1'h0;
endmodule
