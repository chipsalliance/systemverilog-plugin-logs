
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/FunctionScope/dut.sv:1.1-13.10" *)
module dut(clk);
  (* src = "/root/synlig/synlig/tests/simple_tests/FunctionScope/dut.sv:1.19-1.22" *)
  input clk;
  wire clk;
endmodule
