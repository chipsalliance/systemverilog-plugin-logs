
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/NoLatch/dut.sv:1.1-13.10" *)
module dut(clk, a, b);
  (* src = "/root/synlig/synlig/tests/simple_tests/NoLatch/dut.sv:3.17-3.18" *)
  input a;
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/NoLatch/dut.sv:4.17-4.18" *)
  input b;
  wire b;
  (* src = "/root/synlig/synlig/tests/simple_tests/NoLatch/dut.sv:2.17-2.20" *)
  input clk;
  wire clk;
endmodule
