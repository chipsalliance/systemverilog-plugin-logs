
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/DivisionOfSize/top.sv:9.1-13.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/DivisionOfSize/top.sv:9.23-9.24" *)
  output [31:0] o;
  wire [31:0] o;
  (* src = "/root/synlig/synlig/tests/simple_tests/DivisionOfSize/top.sv:11.40-11.58" *)
  wire [2:0] part_buf_data;
  assign o = 32'd7;
  assign part_buf_data = 3'h7;
endmodule
