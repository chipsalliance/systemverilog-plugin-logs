
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypedefWithParameter/top.sv:6.1-9.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefWithParameter/top.sv:6.31-6.32" *)
  output [7:0] o;
  wire [7:0] o;
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefWithParameter/top.sv:7.17-7.26" *)
  (* wiretype = "\\word" *)
  wire [7:0] w;
  assign o = 8'h5c;
  assign w = 8'h5c;
endmodule
