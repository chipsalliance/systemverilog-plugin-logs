
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ArithShiftTernary/top.sv:1.1-7.10" *)
module top(oL, oR);
  (* src = "/root/synlig/synlig/tests/simple_tests/ArithShiftTernary/top.sv:2.14-2.16" *)
  output [31:0] oL;
  wire [31:0] oL;
  (* src = "/root/synlig/synlig/tests/simple_tests/ArithShiftTernary/top.sv:3.14-3.16" *)
  output [31:0] oR;
  wire [31:0] oR;
  assign oL = 32'd512;
  assign oR = 32'd128;
endmodule
