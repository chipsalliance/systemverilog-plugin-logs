
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/HierPathTypespec/dut.sv:33.1-45.10" *)
module dut(clk, i, o);
  (* src = "/root/synlig/synlig/tests/simple_tests/HierPathTypespec/dut.sv:33.24-33.27" *)
  input clk;
  wire clk;
  (* src = "/root/synlig/synlig/tests/simple_tests/HierPathTypespec/dut.sv:33.41-33.42" *)
  input i;
  wire i;
  (* src = "/root/synlig/synlig/tests/simple_tests/HierPathTypespec/dut.sv:33.57-33.58" *)
  output o;
  wire o;
  assign o = i;
endmodule
