
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/Replication/top.sv:1.1-3.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/Replication/top.sv:1.30-1.31" *)
  output [7:0] o;
  wire [7:0] o;
  assign o = 8'h01;
endmodule
