
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/FunctionOnDesignLevel/top.sv:5.1-7.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/FunctionOnDesignLevel/top.sv:5.23-5.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd1;
endmodule
