
(* keep =  1  *)
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:31.1-220.10" *)
module dut();
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:52.45-52.57" *)
  wire [1:0] access_fault;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:44.45-44.59" *)
  wire [33:0] \csr_pmp_addr_i[0] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:44.45-44.59" *)
  wire [33:0] \csr_pmp_addr_i[1] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:44.45-44.59" *)
  wire [33:0] \csr_pmp_addr_i[2] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:44.45-44.59" *)
  wire [33:0] \csr_pmp_addr_i[3] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:43.45-43.58" *)
  (* wiretype = "\\pmp_cfg_t" *)
  wire [23:0] csr_pmp_cfg_i;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:42.45-42.59" *)
  wire [33:0] \pmp_req_addr_i[0] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:42.45-42.59" *)
  wire [33:0] \pmp_req_addr_i[1] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:39.45-39.58" *)
  wire \pmp_req_err_o[0] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:39.45-39.58" *)
  wire \pmp_req_err_o[1] ;
  (* enum_value_00 = "\\PMP_ACC_EXEC" *)
  (* enum_value_01 = "\\PMP_ACC_WRITE" *)
  (* enum_value_10 = "\\PMP_ACC_READ" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:41.45-41.59" *)
  (* wiretype = "\\pmp_req_e" *)
  wire [3:0] pmp_req_type_i;
  (* enum_value_00 = "\\PRIV_LVL_U" *)
  (* enum_value_01 = "\\PRIV_LVL_S" *)
  (* enum_value_10 = "\\PRIV_LVL_H" *)
  (* enum_value_11 = "\\PRIV_LVL_M" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:40.45-40.56" *)
  (* wiretype = "\\priv_lvl_e" *)
  wire [3:0] priv_mode_i;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:46.45-46.61" *)
  wire [33:2] \region_addr_mask[0] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:46.45-46.61" *)
  wire [33:2] \region_addr_mask[1] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:46.45-46.61" *)
  wire [33:2] \region_addr_mask[2] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:46.45-46.61" *)
  wire [33:2] \region_addr_mask[3] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:50.45-50.61" *)
  wire [7:0] region_match_all;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:49.45-49.60" *)
  wire [7:0] region_match_eq;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:47.45-47.60" *)
  wire [7:0] region_match_gt;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:48.45-48.60" *)
  wire [7:0] region_match_lt;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:51.45-51.62" *)
  wire [7:0] region_perm_check;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:45.45-45.62" *)
  wire [33:0] \region_start_addr[0] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:45.45-45.62" *)
  wire [33:0] \region_start_addr[1] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:45.45-45.62" *)
  wire [33:0] \region_start_addr[2] ;
  (* src = "/root/synlig/synlig/tests/simple_tests/hier_path/dut.sv:45.45-45.62" *)
  wire [33:0] \region_start_addr[3] ;
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  assign access_fault = 2'h0;
  assign \csr_pmp_addr_i[0]  = 34'h000000000;
  assign \csr_pmp_addr_i[1]  = 34'h111111111;
  assign \csr_pmp_addr_i[2]  = 34'h111111111;
  assign \csr_pmp_addr_i[3]  = 34'h111111111;
  assign csr_pmp_cfg_i = 24'hbffdc8;
  assign \pmp_req_addr_i[0]  = 34'h000000000;
  assign \pmp_req_addr_i[1]  = 34'h111111111;
  assign \pmp_req_err_o[0]  = 1'h0;
  assign \pmp_req_err_o[1]  = 1'h0;
  assign pmp_req_type_i = 4'h0;
  assign priv_mode_i = 4'hb;
  assign \region_addr_mask[0]  = 32'd4294967295;
  assign \region_addr_mask[1]  = 32'd4294967295;
  assign \region_addr_mask[2]  = 32'd4294967294;
  assign \region_addr_mask[3]  = 32'd4294967295;
  assign region_match_all = 8'h60;
  assign region_match_eq = 8'he1;
  assign region_match_gt = 8'h10;
  assign region_match_lt = 8'h0e;
  assign region_perm_check = 8'hee;
  assign \region_start_addr[0]  = 34'h000000000;
  assign \region_start_addr[1]  = 34'h111111111;
  assign \region_start_addr[2]  = 34'h111111111;
  assign \region_start_addr[3]  = 34'h111111111;
endmodule
