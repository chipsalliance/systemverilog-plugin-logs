
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TaskImportDPI/top.sv:1.1-7.10" *)
module top(a);
  (* src = "/root/synlig/synlig/tests/simple_tests/TaskImportDPI/top.sv:1.23-1.24" *)
  output [31:0] a;
  wire [31:0] a;
  (* nosync = 32'd1 *)
  (* src = "/root/synlig/synlig/tests/simple_tests/TaskImportDPI/top.sv:2.56-2.57" *)
  wire [31:0] \test_output_argument$func$/root/synlig/synlig/tests/simple_tests/TaskImportDPI/top.sv:5$1.o ;
  assign \test_output_argument$func$/root/synlig/synlig/tests/simple_tests/TaskImportDPI/top.sv:5$1.o  = a;
endmodule
