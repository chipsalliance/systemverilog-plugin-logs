
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/Shortint/top.sv:1.1-3.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/Shortint/top.sv:1.28-1.29" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd1;
endmodule
