
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/onenet/top.sv:1.1-3.10" *)
module top(a, b);
  (* src = "/root/synlig/synlig/tests/simple_tests/onenet/top.sv:1.18-1.19" *)
  input a;
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/onenet/top.sv:1.28-1.29" *)
  output b;
  wire b;
  assign b = a;
endmodule
