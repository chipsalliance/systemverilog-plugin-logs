
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ParameterInitializedByPartSelectOfParameters/top.sv:1.1-6.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterInitializedByPartSelectOfParameters/top.sv:1.31-1.32" *)
  output [5:0] o;
  wire [5:0] o;
  assign o = 6'h14;
endmodule
