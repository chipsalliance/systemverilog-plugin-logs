
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/Shortreal/top.sv:1.1-4.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/Shortreal/top.sv:2.14-2.21" *)
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/Shortreal/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign a = 1'h1;
  assign o = 32'd2;
endmodule
