
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/GetC/top.sv:1.1-4.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/GetC/top.sv:2.11-2.21" *)
  wire [31:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/GetC/top.sv:1.24-1.25" *)
  output [7:0] o;
  wire [7:0] o;
  assign a = 32'd1415934836;
  assign o = 8'h74;
endmodule
