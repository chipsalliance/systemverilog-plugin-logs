
(* cells_not_processed =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/UnionInPackageWithMultirange/top.sv:34.1-36.10" *)
module top(b, a);
  (* src = "/root/synlig/synlig/tests/simple_tests/UnionInPackageWithMultirange/top.sv:34.35-34.36" *)
  (* wiretype = "\\top_flag_t" *)
  input [95:0] a;
  wire [95:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/UnionInPackageWithMultirange/top.sv:34.63-34.64" *)
  (* wiretype = "\\top_flag_t" *)
  output [95:0] b;
  wire [95:0] b;
  assign b = a;
endmodule
