
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ImportedParameter/top.sv:5.1-8.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ImportedParameter/top.sv:5.23-5.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd4;
endmodule
