
(* keep =  1  *)
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ParameterUnpackedLogicArray/top.sv:1.1-22.10" *)
module top(a, b, c, d);
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterUnpackedLogicArray/top.sv:1.25-1.26" *)
  output a;
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterUnpackedLogicArray/top.sv:1.28-1.29" *)
  output b;
  wire b;
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterUnpackedLogicArray/top.sv:1.31-1.32" *)
  output c;
  wire c;
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterUnpackedLogicArray/top.sv:1.34-1.35" *)
  output d;
  wire d;
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  always @*
    if (1'h1) begin
      assert (1'h1);
    end
  assign a = 1'h1;
  assign b = 1'h0;
  assign c = 1'h0;
  assign d = 1'h0;
endmodule
