
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/UnitForLoop/dut.v:1.1-17.10" *)
module dut(a, b);
  (* src = "/root/synlig/synlig/tests/simple_tests/UnitForLoop/dut.v:1.18-1.19" *)
  input a;
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/UnitForLoop/dut.v:1.28-1.29" *)
  output b;
  wire b;
  assign b = a;
endmodule
