
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/DisplayWithHexFormatSpecifier/top.sv:1.1-5.10" *)
module top();
endmodule
