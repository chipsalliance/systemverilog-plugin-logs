
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/conditional_if_else/if_else.sv:6.1-13.10" *)
module top();
  (* src = "/root/synlig/synlig/tests/simple_tests/conditional_if_else/if_else.sv:7.7-7.8" *)
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/conditional_if_else/if_else.sv:8.6-8.11" *)
  wire b;
  assign a = 1'h1;
  assign b = 1'h1;
endmodule
