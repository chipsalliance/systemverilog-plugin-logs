
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ParameterConditionalAssignment/top.sv:1.1-11.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterConditionalAssignment/top.sv:4.17-4.18" *)
  output o;
  wire o;
  assign o = 1'h1;
endmodule
