
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ParameterOfSizeOfParametrizedPort/top.sv:1.1-8.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterOfSizeOfParametrizedPort/top.sv:4.25-4.26" *)
  output [14:0] o;
  wire [14:0] o;
  assign o = 15'h7fff;
endmodule
