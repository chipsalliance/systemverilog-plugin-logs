
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CastSize/top.sv:1.1-6.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CastSize/top.sv:2.17-2.27" *)
  wire [15:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/CastSize/top.sv:1.31-1.32" *)
  output [4:0] o;
  wire [4:0] o;
  assign a = 16'h00ab;
  assign o = 5'h0b;
endmodule
