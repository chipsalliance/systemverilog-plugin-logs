
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/AssignmentPattern/top.sv:1.1-24.10" *)
module top(b);
  (* src = "/root/synlig/synlig/tests/simple_tests/AssignmentPattern/top.sv:9.14-9.15" *)
  (* wiretype = "\\struct_t" *)
  wire [3:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/AssignmentPattern/top.sv:1.25-1.26" *)
  output [3:0] b;
  wire [3:0] b;
  assign a = 4'h5;
  assign b = 4'h5;
endmodule
