
(* dynports =  1  *)
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/StreamOp/dut.sv:1.1-16.10" *)
module dut(a, b, c, d);
  (* src = "/root/synlig/synlig/tests/simple_tests/StreamOp/dut.sv:1.32-1.33" *)
  output [31:0] a;
  wire [31:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/StreamOp/dut.sv:1.35-1.36" *)
  output [31:0] b;
  wire [31:0] b;
  (* src = "/root/synlig/synlig/tests/simple_tests/StreamOp/dut.sv:1.58-1.59" *)
  output [63:0] c;
  wire [63:0] c;
  (* src = "/root/synlig/synlig/tests/simple_tests/StreamOp/dut.sv:1.61-1.62" *)
  output [63:0] d;
  wire [63:0] d;
  (* src = "/root/synlig/synlig/tests/simple_tests/StreamOp/dut.sv:2.15-2.16" *)
  wire [31:0] x;
  (* src = "/root/synlig/synlig/tests/simple_tests/StreamOp/dut.sv:3.15-3.16" *)
  wire [31:0] y;
  assign a = 32'd4286523927;
  assign b = 32'd388661247;
  assign c = 64'h172a7fffff7f2a17;
  assign d = 64'h172a7fffff7f2a17;
  assign x = 32'd388661247;
  assign y = 32'd4286523927;
endmodule
