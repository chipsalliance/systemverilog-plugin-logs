
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ParameterInitializationWithNegation/top.sv:1.1-4.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ParameterInitializationWithNegation/top.sv:1.32-1.33" *)
  output [17:0] o;
  wire [17:0] o;
  assign o = 18'h3fff0;
endmodule
