
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/conditional_if/if.sv:6.1-12.10" *)
module top();
  (* src = "/root/synlig/synlig/tests/simple_tests/conditional_if/if.sv:7.10-7.11" *)
  wire a;
  (* init = 1'h0 *)
  (* src = "/root/synlig/synlig/tests/simple_tests/conditional_if/if.sv:8.9-8.14" *)
  (* unused_bits = "0" *)
  wire b;
  assign a = 1'h0;
endmodule
