
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CastInFunctionToParameterWidth/top.sv:1.1-12.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CastInFunctionToParameterWidth/top.sv:5.33-5.34" *)
  output [14:0] o;
  wire [14:0] o;
  assign o = 15'h0003;
endmodule
