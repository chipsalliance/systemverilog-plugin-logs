
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/IndexedPartSelectOfArrayElement/top.sv:1.1-8.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/IndexedPartSelectOfArrayElement/top.sv:6.13-6.14" *)
  (* wiretype = "\\tl_h2d_t" *)
  wire [15:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/IndexedPartSelectOfArrayElement/top.sv:1.31-1.32" *)
  output [1:0] o;
  wire [1:0] o;
  assign a = 16'h0012;
  assign o = 2'h0;
endmodule
