
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/OneSysFunc/dut.v:1.1-3.10" *)
module dut(a, b);
  (* src = "/root/synlig/synlig/tests/simple_tests/OneSysFunc/dut.v:1.19-1.20" *)
  input a;
  wire a;
  (* src = "/root/synlig/synlig/tests/simple_tests/OneSysFunc/dut.v:1.29-1.30" *)
  output b;
  wire b;
  assign b = a;
endmodule
