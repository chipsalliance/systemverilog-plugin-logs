
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumConstX/top.sv:1.1-15.10" *)
module top(clk, out);
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumConstX/top.sv:1.24-1.27" *)
  input clk;
  wire clk;
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumConstX/top.sv:1.47-1.50" *)
  output [3:0] out;
  wire [3:0] out;
  assign out = 4'b1xxx;
endmodule
