
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/TypedefedFunctionArgument/top.sv:1.1-9.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefedFunctionArgument/top.sv:7.9-7.10" *)
  (* wiretype = "\\word" *)
  wire [31:0] a;
  (* nosync = 32'd1 *)
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefedFunctionArgument/top.sv:3.54-3.55" *)
  (* wiretype = "\\word" *)
  wire [31:0] \check_if_abcd$func$/root/synlig/synlig/tests/simple_tests/TypedefedFunctionArgument/top.sv:8$2.x ;
  (* src = "/root/synlig/synlig/tests/simple_tests/TypedefedFunctionArgument/top.sv:1.25-1.26" *)
  output o;
  wire o;
  assign a = 32'd43981;
  assign \check_if_abcd$func$/root/synlig/synlig/tests/simple_tests/TypedefedFunctionArgument/top.sv:8$2.x  = 32'hxxxxxxxx;
  assign o = 1'h1;
endmodule
