
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/FunctionWithoutReturn/top.sv:7.1-9.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/FunctionWithoutReturn/top.sv:7.19-7.20" *)
  output o;
  wire o;
  assign o = 1'h1;
endmodule
