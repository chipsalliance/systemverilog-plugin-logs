
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/AssignArraySelPlus/top.sv:1.1-6.10" *)
module top(data);
  (* src = "/root/synlig/synlig/tests/simple_tests/AssignArraySelPlus/top.sv:1.32-1.36" *)
  output [63:0] data;
  wire [63:0] data;
  assign data[43:40] = 4'hf;
endmodule
