
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/EnumArrayListedElements/top.sv:8.1-11.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumArrayListedElements/top.sv:8.23-8.24" *)
  output [31:0] o;
  wire [31:0] o;
  (* enum_value_1010 = "\\On" *)
  (* enum_value_1111 = "\\Off" *)
  (* src = "/root/synlig/synlig/tests/simple_tests/EnumArrayListedElements/top.sv:9.26-9.56" *)
  (* wiretype = "\\lc_tx_t" *)
  wire [7:0] x;
  assign o = 32'd175;
  assign x = 8'haf;
endmodule
