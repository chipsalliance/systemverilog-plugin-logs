
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/CaseWithGeneratedWire/top.sv:1.1-15.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/CaseWithGeneratedWire/top.sv:5.21-5.22" *)
  wire \gen_blk[0].z ;
  (* src = "/root/synlig/synlig/tests/simple_tests/CaseWithGeneratedWire/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign \gen_blk[0].z  = 1'h1;
  assign o = 32'd1;
endmodule
