
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ImportedDoubleCastedParameter/top.sv:11.1-14.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ImportedDoubleCastedParameter/top.sv:11.23-11.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign o = 32'd1073807361;
endmodule
