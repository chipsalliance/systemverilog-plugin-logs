
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/AssignBitSelectPartSelect/top.sv:1.1-4.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/AssignBitSelectPartSelect/top.sv:1.30-1.31" *)
  output [1:0] o;
  wire [1:0] o;
  (* src = "/root/synlig/synlig/tests/simple_tests/AssignBitSelectPartSelect/top.sv:2.21-2.27" *)
  wire [9:0] x;
  assign o = 2'h3;
  assign x = 10'h3ff;
endmodule
