
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ReturnFunctionCall/top.sv:11.1-13.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ReturnFunctionCall/top.sv:11.25-11.26" *)
  output o;
  wire o;
  assign o = 1'h1;
endmodule
