
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/ForkJoinTypes/top.sv:1.1-14.10" *)
module top(o);
  (* src = "/root/synlig/synlig/tests/simple_tests/ForkJoinTypes/top.sv:2.8-2.9" *)
  wire [31:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/ForkJoinTypes/top.sv:1.23-1.24" *)
  output [31:0] o;
  wire [31:0] o;
  assign a = 32'd0;
  assign o = 32'd0;
endmodule
