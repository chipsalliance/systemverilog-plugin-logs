
(* top =  1  *)
(* src = "/root/synlig/synlig/tests/simple_tests/IndexedPartSelect/top.sv:1.1-6.10" *)
module top(b, c);
  (* src = "/root/synlig/synlig/tests/simple_tests/IndexedPartSelect/top.sv:2.14-2.15" *)
  wire [7:0] a;
  (* src = "/root/synlig/synlig/tests/simple_tests/IndexedPartSelect/top.sv:1.25-1.26" *)
  output [3:0] b;
  wire [3:0] b;
  (* src = "/root/synlig/synlig/tests/simple_tests/IndexedPartSelect/top.sv:1.41-1.42" *)
  output [3:0] c;
  wire [3:0] c;
  assign a = 8'h0f;
  assign b = 4'h3;
  assign c = 4'h3;
endmodule
